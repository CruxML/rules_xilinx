module empty_top ();

endmodule

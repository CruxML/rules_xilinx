module zcu111_submodule (
    input  logic a,
    output logic b
);

  assign b = !a;

endmodule

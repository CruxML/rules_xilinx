module empty_top (
    output logic [7:0] leds
);

  assign leds = 8'hA5;

endmodule
